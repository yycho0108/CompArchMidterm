`ifndef __ENCODER_V__
`define __ENCODER_V__
`include "defs.v"

// 0001 --> 00
// 0010 --> 01, etc.

module encoder
(

);

endmodule
`endif
