`include "defs.v"

// 0001 --> 00
// 0010 --> 01, etc.

module encoder
(

);

endmodule
